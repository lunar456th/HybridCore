module CLA(n, z, o, a, b);
	input [3:0] a, b;
	input o;
	wire [3:0] p, g, c;
	wire [9:0] m;
	output [3:0] n;
	output z;
	xor (p[0], a[0], b[0]);
	and (g[0], a[0], b[0]);
	xor (p[1], a[1], b[1]);
	and (g[1], a[1], b[1]);
	xor (p[2], a[2], b[2]);
	and (g[2], a[2], b[2]);
	xor (p[3], a[3], b[3]);
	and (g[3], a[3], b[3]);
	and (m[0], o, p[0]);
	or (c[0], m[0], g[0]);
	and (m[1], g[0], p[1]);
	and (m[2], o, p[0], p[1]);
	or (c[1], g[1], m[1], m[2]);
	and (m[3], g[1], p[2]);
	and (m[4], g[0], p[1], p[2]);
	and (m[5], o, p[1], p[2], p[0]);
	or (c[2], g[2], m[3], m[4], m[5]);
	and (m[6], g[2], p[3]);
	and (m[7], g[1], p[2], p[3]);
	and (m[8], g[0], p[1], p[2], p[3]);
	and (m[9], o, p[0], p[1], p[2], p[3]);
	or (c[3], g[3], m[6], m[7], m[8], m[9]);
	xor (n[0], p[0], o);
	xor (n[1], p[1], c[0]);
	xor (n[2], p[2], c[1]);
	xor (n[3], p[3], c[2]);
	assign z = c[3];
endmodule