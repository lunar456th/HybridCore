/*
	Name		:	Divider
	File		:	divider.v
	Word size	:	16-bit
	Algorithm	:	Look-up table
	Url			:	https://github.com/srichandra/fast-division
*/

module divider (
	input wire clk;
	input wire en;
	input wire [15:0] a;
	input wire [15:0] b;
	output wire [31:0] xyout;
    );
	
	reg [31:0] xyouti;
	reg [15:0] out;
	wire [31:0] temp;
	
	mult mult(out, a, temp);
	
	always @ (b)
	begin
		casex(b)
			16'b0000000000000010: out <= 16'h8000;
			16'b0000000000000011: out <= 16'h5555;
			16'b0000000000000100: out <= 16'h4000;
			16'b0000000000000101: out <= 16'h3333;
			16'b0000000000000110: out <= 16'h2AAA;
			16'b0000000000000111: out <= 16'h2492;
			16'b0000000000001000: out <= 16'h2000;
			16'b0000000000001001: out <= 16'h1C71;
			16'b0000000000001010: out <= 16'h1999;
			16'b0000000000001011: out <= 16'h1745;
			16'b0000000000001100: out <= 16'h1555;
			16'b0000000000001101: out <= 16'h13B1;
			16'b0000000000001110: out <= 16'h1249;
			16'b0000000000001111: out <= 16'h1111;
			16'b0000000000010000: out <= 16'h1000;
			16'b0000000000010001: out <= 16'h0F0F;
			16'b0000000000010010: out <= 16'h0E38;
			16'b0000000000010011: out <= 16'h0D79;
			16'b0000000000010100: out <= 16'h0CCC;
			16'b0000000000010101: out <= 16'h0C30;
			16'b0000000000010110: out <= 16'h0BA2;
			16'b0000000000010111: out <= 16'h0B21;
			16'b0000000000011000: out <= 16'h0AAA;
			16'b0000000000011001: out <= 16'h0A3D;
			16'b0000000000011010: out <= 16'h09D8;
			16'b0000000000011011: out <= 16'h097B;
			16'b0000000000011100: out <= 16'h0924;
			16'b0000000000011101: out <= 16'h08D3;
			16'b0000000000011110: out <= 16'h0888;
			16'b0000000000011111: out <= 16'h0842;
			16'b0000000000100000: out <= 16'h0800;
			16'b0000000000100001: out <= 16'h07C1;
			16'b0000000000100010: out <= 16'h0787;
			16'b0000000000100011: out <= 16'h0750;
			16'b0000000000100100: out <= 16'h071C;
			16'b0000000000100101: out <= 16'h06EB;
			16'b0000000000100110: out <= 16'h06BC;
			16'b0000000000100111: out <= 16'h0690;
			16'b0000000000101000: out <= 16'h0666;
			16'b0000000000101001: out <= 16'h063E;
			16'b0000000000101010: out <= 16'h0618;
			16'b0000000000101011: out <= 16'h05F4;
			16'b0000000000101100: out <= 16'h05D1;
			16'b0000000000101101: out <= 16'h05B0;
			16'b0000000000101110: out <= 16'h0590;
			16'b0000000000101111: out <= 16'h0572;
			16'b0000000000110000: out <= 16'h0555;
			16'b0000000000110001: out <= 16'h0539;
			16'b0000000000110010: out <= 16'h051E;
			16'b0000000000110011: out <= 16'h0505;
			16'b0000000000110100: out <= 16'h04EC;
			16'b0000000000110101: out <= 16'h04D4;
			16'b0000000000110110: out <= 16'h04BD;
			16'b0000000000110111: out <= 16'h04A7;
			16'b0000000000111000: out <= 16'h0492;
			16'b0000000000111001: out <= 16'h047D;
			16'b0000000000111010: out <= 16'h0469;
			16'b0000000000111011: out <= 16'h0456;
			16'b0000000000111100: out <= 16'h0444;
			16'b0000000000111101: out <= 16'h0432;
			16'b0000000000111110: out <= 16'h0421;
			16'b0000000000111111: out <= 16'h0410;
			16'b0000000001000000: out <= 16'h0400;
			16'b0000000001000001: out <= 16'h03F0;
			16'b0000000001000010: out <= 16'h03E0;
			16'b0000000001000011: out <= 16'h03D2;
			16'b0000000001000100: out <= 16'h03C3;
			16'b0000000001000101: out <= 16'h03B5;
			16'b0000000001000110: out <= 16'h03A8;
			16'b0000000001000111: out <= 16'h039B;
			16'b0000000001001000: out <= 16'h038E;
			16'b0000000001001001: out <= 16'h0381;
			16'b0000000001001010: out <= 16'h0375;
			16'b0000000001001011: out <= 16'h0369;
			16'b0000000001001100: out <= 16'h035E;
			16'b0000000001001101: out <= 16'h0353;
			16'b0000000001001110: out <= 16'h0348;
			16'b0000000001001111: out <= 16'h033D;
			16'b0000000001010000: out <= 16'h0333;
			16'b0000000001010001: out <= 16'h0329;
			16'b0000000001010010: out <= 16'h031F;
			16'b0000000001010011: out <= 16'h0315;
			16'b0000000001010100: out <= 16'h030C;
			16'b0000000001010101: out <= 16'h0303;
			16'b0000000001010110: out <= 16'h02FA;
			16'b0000000001010111: out <= 16'h02F1;
			16'b0000000001011000: out <= 16'h02E8;
			16'b0000000001011001: out <= 16'h02E0;
			16'b0000000001011010: out <= 16'h02D8;
			16'b0000000001011011: out <= 16'h02D0;
			16'b0000000001011100: out <= 16'h02C8;
			16'b0000000001011101: out <= 16'h02C0;
			16'b0000000001011110: out <= 16'h02B9;
			16'b0000000001011111: out <= 16'h02B1;
			16'b0000000001100000: out <= 16'h02AA;
			16'b0000000001100001: out <= 16'h02A3;
			16'b0000000001100010: out <= 16'h029C;
			16'b0000000001100011: out <= 16'h0295;
			16'b0000000001100100: out <= 16'h028F;
			16'b0000000001100101: out <= 16'h0288;
			16'b0000000001100110: out <= 16'h0282;
			16'b0000000001100111: out <= 16'h027C;
			16'b0000000001101000: out <= 16'h0276;
			16'b0000000001101001: out <= 16'h0270;
			16'b0000000001101010: out <= 16'h026A;
			16'b0000000001101011: out <= 16'h0264;
			16'b0000000001101100: out <= 16'h025E;
			16'b0000000001101101: out <= 16'h0259;
			16'b0000000001101110: out <= 16'h0253;
			16'b0000000001101111: out <= 16'h024E;
			16'b0000000001110000: out <= 16'h0249;
			16'b0000000001110001: out <= 16'h0243;
			16'b0000000001110010: out <= 16'h023E;
			16'b0000000001110011: out <= 16'h0239;
			16'b0000000001110100: out <= 16'h0234;
			16'b0000000001110101: out <= 16'h0230;
			16'b0000000001110110: out <= 16'h022B;
			16'b0000000001110111: out <= 16'h0226;
			16'b0000000001111000: out <= 16'h0222;
			16'b0000000001111001: out <= 16'h021D;
			16'b0000000001111010: out <= 16'h0219;
			16'b0000000001111011: out <= 16'h0214;
			16'b0000000001111100: out <= 16'h0210;
			16'b0000000001111101: out <= 16'h020C;
			16'b0000000001111110: out <= 16'h0208;
			16'b0000000001111111: out <= 16'h0204;
			16'b0000000010000000: out <= 16'h0200;
			16'b0000000010000001: out <= 16'h01FC;
			16'b0000000010000010: out <= 16'h01F8;
			16'b0000000010000011: out <= 16'h01F4;
			16'b0000000010000100: out <= 16'h01F0;
			16'b0000000010000101: out <= 16'h01EC;
			16'b0000000010000110: out <= 16'h01E9;
			16'b0000000010000111: out <= 16'h01E5;
			16'b0000000010001000: out <= 16'h01E1;
			16'b0000000010001001: out <= 16'h01DE;
			16'b0000000010001010: out <= 16'h01DA;
			16'b0000000010001011: out <= 16'h01D7;
			16'b0000000010001100: out <= 16'h01D4;
			16'b0000000010001101: out <= 16'h01D0;
			16'b0000000010001110: out <= 16'h01CD;
			16'b0000000010001111: out <= 16'h01CA;
			16'b0000000010010000: out <= 16'h01C7;
			16'b0000000010010001: out <= 16'h01C3;
			16'b0000000010010010: out <= 16'h01C0;
			16'b0000000010010011: out <= 16'h01BD;
			16'b0000000010010100: out <= 16'h01BA;
			16'b0000000010010101: out <= 16'h01B7;
			16'b0000000010010110: out <= 16'h01B4;
			16'b0000000010010111: out <= 16'h01B2;
			16'b0000000010011000: out <= 16'h01AF;
			16'b0000000010011001: out <= 16'h01AC;
			16'b0000000010011010: out <= 16'h01A9;
			16'b0000000010011011: out <= 16'h01A6;
			16'b0000000010011100: out <= 16'h01A4;
			16'b0000000010011101: out <= 16'h01A1;
			16'b0000000010011110: out <= 16'h019E;
			16'b0000000010011111: out <= 16'h019C;
			16'b0000000010100000: out <= 16'h0199;
			16'b0000000010100001: out <= 16'h0197;
			16'b0000000010100010: out <= 16'h0194;
			16'b0000000010100011: out <= 16'h0192;
			16'b0000000010100100: out <= 16'h018F;
			16'b0000000010100101: out <= 16'h018D;
			16'b0000000010100110: out <= 16'h018A;
			16'b0000000010100111: out <= 16'h0188;
			16'b0000000010101000: out <= 16'h0186;
			16'b0000000010101001: out <= 16'h0183;
			16'b0000000010101010: out <= 16'h0181;
			16'b0000000010101011: out <= 16'h017F;
			16'b0000000010101100: out <= 16'h017D;
			16'b0000000010101101: out <= 16'h017A;
			16'b0000000010101110: out <= 16'h0178;
			16'b0000000010101111: out <= 16'h0176;
			16'b0000000010110000: out <= 16'h0174;
			16'b0000000010110001: out <= 16'h0172;
			16'b0000000010110010: out <= 16'h0170;
			16'b0000000010110011: out <= 16'h016E;
			16'b0000000010110100: out <= 16'h016C;
			16'b0000000010110101: out <= 16'h016A;
			16'b0000000010110110: out <= 16'h0168;
			16'b0000000010110111: out <= 16'h0166;
			16'b0000000010111000: out <= 16'h0164;
			16'b0000000010111001: out <= 16'h0162;
			16'b0000000010111010: out <= 16'h0160;
			16'b0000000010111011: out <= 16'h015E;
			16'b0000000010111100: out <= 16'h015C;
			16'b0000000010111101: out <= 16'h015A;
			16'b0000000010111110: out <= 16'h0158;
			16'b0000000010111111: out <= 16'h0157;
			16'b0000000011000000: out <= 16'h0155;
			16'b0000000011000001: out <= 16'h0153;
			16'b0000000011000010: out <= 16'h0151;
			16'b0000000011000011: out <= 16'h0150;
			16'b0000000011000100: out <= 16'h014E;
			16'b0000000011000101: out <= 16'h014C;
			16'b0000000011000110: out <= 16'h014A;
			16'b0000000011000111: out <= 16'h0149;
			16'b0000000011001000: out <= 16'h0147;
			16'b0000000011001001: out <= 16'h0146;
			16'b0000000011001010: out <= 16'h0144;
			16'b0000000011001011: out <= 16'h0142;
			16'b0000000011001100: out <= 16'h0141;
			16'b0000000011001101: out <= 16'h013F;
			16'b0000000011001110: out <= 16'h013E;
			16'b0000000011001111: out <= 16'h013C;
			16'b0000000011010000: out <= 16'h013B;
			16'b0000000011010001: out <= 16'h0139;
			16'b0000000011010010: out <= 16'h0138;
			16'b0000000011010011: out <= 16'h0136;
			16'b0000000011010100: out <= 16'h0135;
			16'b0000000011010101: out <= 16'h0133;
			16'b0000000011010110: out <= 16'h0132;
			16'b0000000011010111: out <= 16'h0130;
			16'b0000000011011000: out <= 16'h012F;
			16'b0000000011011001: out <= 16'h012E;
			16'b0000000011011010: out <= 16'h012C;
			16'b0000000011011011: out <= 16'h012B;
			16'b0000000011011100: out <= 16'h0129;
			16'b0000000011011101: out <= 16'h0128;
			16'b0000000011011110: out <= 16'h0127;
			16'b0000000011011111: out <= 16'h0125;
			16'b0000000011100000: out <= 16'h0124;
			16'b0000000011100001: out <= 16'h0123;
			16'b0000000011100010: out <= 16'h0121;
			16'b0000000011100011: out <= 16'h0120;
			16'b0000000011100100: out <= 16'h011F;
			16'b0000000011100101: out <= 16'h011E;
			16'b0000000011100110: out <= 16'h011C;
			16'b0000000011100111: out <= 16'h011B;
			16'b0000000011101000: out <= 16'h011A;
			16'b0000000011101001: out <= 16'h0119;
			16'b0000000011101010: out <= 16'h0118;
			16'b0000000011101011: out <= 16'h0116;
			16'b0000000011101100: out <= 16'h0115;
			16'b0000000011101101: out <= 16'h0114;
			16'b0000000011101110: out <= 16'h0113;
			16'b0000000011101111: out <= 16'h0112;
			16'b0000000011110000: out <= 16'h0111;
			16'b0000000011110001: out <= 16'h010F;
			16'b0000000011110010: out <= 16'h010E;
			16'b0000000011110011: out <= 16'h010D;
			16'b0000000011110100: out <= 16'h010C;
			16'b0000000011110101: out <= 16'h010B;
			16'b0000000011110110: out <= 16'h010A;
			16'b0000000011110111: out <= 16'h0109;
			16'b0000000011111000: out <= 16'h0108;
			16'b0000000011111001: out <= 16'h0107;
			16'b0000000011111010: out <= 16'h0106;
			16'b0000000011111011: out <= 16'h0105;
			16'b0000000011111100: out <= 16'h0104;
			16'b0000000011111101: out <= 16'h0103;
			16'b0000000011111110: out <= 16'h0102;
			16'b0000000011111111: out <= 16'h0101;
			16'b0000000100000000: out <= 16'h0100;
			16'b0000000100000001: out <= 16'h00FF;
			16'b0000000100000010: out <= 16'h00FE;
			16'b0000000100000011: out <= 16'h00FD;
			16'b0000000100000100: out <= 16'h00FC;
			16'b0000000100000101: out <= 16'h00FB;
			16'b0000000100000110: out <= 16'h00FA;
			16'b0000000100000111: out <= 16'h00F9;
			16'b0000000100001000: out <= 16'h00F8;
			16'b0000000100001001: out <= 16'h00F7;
			16'b0000000100001010: out <= 16'h00F6;
			16'b0000000100001011: out <= 16'h00F5;
			16'b0000000100001100: out <= 16'h00F4;
			16'b0000000100001101: out <= 16'h00F3;
			16'b0000000100001110: out <= 16'h00F2;
			16'b0000000100001111: out <= 16'h00F1;
			16'b000000010001000x: out <= 16'h00F0;
			16'b0000000100010010: out <= 16'h00EF;
			16'b0000000100010011: out <= 16'h00EE;
			16'b0000000100010100: out <= 16'h00ED;
			16'b0000000100010101: out <= 16'h00EC;
			16'b0000000100010110: out <= 16'h00EB;
			16'b000000010001011x: out <= 16'h00EA;
			16'b0000000100011001: out <= 16'h00E9;
			16'b0000000100011010: out <= 16'h00E8;
			16'b0000000100011011: out <= 16'h00E7;
			16'b0000000100011100: out <= 16'h00E6;
			16'b0000000100011101: out <= 16'h00E5;
			16'b0000000100011110: out <= 16'h00E5;
			16'b0000000100011111: out <= 16'h00E4;
			16'b0000000100100000: out <= 16'h00E3;
			16'b0000000100100001: out <= 16'h00E2;
			16'b000000010010001x: out <= 16'h00E1;
			16'b0000000100100100: out <= 16'h00E0;
			16'b0000000100100101: out <= 16'h00DF;
			16'b000000010010011x: out <= 16'h00DE;
			16'b0000000100101000: out <= 16'h00DD;
			16'b0000000100101001: out <= 16'h00DC;
			16'b000000010010101x: out <= 16'h00DB;
			16'b0000000100101100: out <= 16'h00DA;
			16'b0000000100101101: out <= 16'h00D9;
			16'b0000000100101110: out <= 16'h00D9;
			16'b0000000100101111: out <= 16'h00D8;
			16'b0000000100110000: out <= 16'h00D7;
			16'b0000000100110001: out <= 16'h00D6;
			16'b0000000100110010: out <= 16'h00D6;
			16'b0000000100110011: out <= 16'h00D5;
			16'b000000010011010x: out <= 16'h00D4;
			16'b0000000100110110: out <= 16'h00D3;
			16'b0000000100110111: out <= 16'h00D2;
			16'b0000000100111000: out <= 16'h00D2;
			16'b0000000100111001: out <= 16'h00D1;
			16'b000000010011101x: out <= 16'h00D0;
			16'b0000000100111100: out <= 16'h00CF;
			16'b0000000100111101: out <= 16'h00CE;
			16'b0000000100111110: out <= 16'h00CE;
			16'b0000000100111111: out <= 16'h00CD;
			16'b000000010100000x: out <= 16'h00CC;
			16'b0000000101000010: out <= 16'h00CB;
			16'b0000000101000011: out <= 16'h00CA;
			16'b0000000101000100: out <= 16'h00CA;
			16'b0000000101000101: out <= 16'h00C9;
			16'b0000000101000110: out <= 16'h00C9;
			16'b0000000101000111: out <= 16'h00C8;
			16'b000000010100100x: out <= 16'h00C7;
			16'b0000000101001010: out <= 16'h00C6;
			16'b0000000101001011: out <= 16'h00C5;
			16'b0000000101001100: out <= 16'h00C5;
			16'b0000000101001101: out <= 16'h00C4;
			16'b0000000101001110: out <= 16'h00C4;
			16'b0000000101001111: out <= 16'h00C3;
			16'b0000000101010000: out <= 16'h00C3;
			16'b0000000101010001: out <= 16'h00C2;
			16'b000000010101001x: out <= 16'h00C1;
			16'b000000010101010x: out <= 16'h00C0;
			16'b000000010101011x: out <= 16'h00BF;
			16'b0000000101011000: out <= 16'h00BE;
			16'b0000000101011001: out <= 16'h00BD;
			16'b0000000101011010: out <= 16'h00BD;
			16'b0000000101011011: out <= 16'h00BC;
			16'b0000000101011100: out <= 16'h00BC;
			16'b0000000101011101: out <= 16'h00BB;
			16'b0000000101011110: out <= 16'h00BB;
			16'b0000000101011111: out <= 16'h00BA;
			16'b0000000101100000: out <= 16'h00BA;
			16'b0000000101100001: out <= 16'h00B9;
			16'b0000000101100010: out <= 16'h00B9;
			16'b0000000101100011: out <= 16'h00B8;
			16'b0000000101100100: out <= 16'h00B8;
			16'b0000000101100101: out <= 16'h00B7;
			16'b0000000101100110: out <= 16'h00B7;
			16'b0000000101100111: out <= 16'h00B6;
			16'b0000000101101000: out <= 16'h00B6;
			16'b0000000101101001: out <= 16'h00B5;
			16'b0000000101101010: out <= 16'h00B5;
			16'b0000000101101011: out <= 16'h00B4;
			16'b0000000101101100: out <= 16'h00B4;
			16'b0000000101101101: out <= 16'h00B3;
			16'b0000000101101110: out <= 16'h00B3;
			16'b0000000101101111: out <= 16'h00B2;
			16'b0000000101110000: out <= 16'h00B2;
			16'b0000000101110001: out <= 16'h00B1;
			16'b0000000101110010: out <= 16'h00B1;
			16'b0000000101110011: out <= 16'h00B0;
			16'b0000000101110100: out <= 16'h00B0;
			16'b0000000101110101: out <= 16'h00AF;
			16'b0000000101110110: out <= 16'h00AF;
			16'b0000000101110111: out <= 16'h00AE;
			16'b0000000101111000: out <= 16'h00AE;
			16'b0000000101111001: out <= 16'h00AD;
			16'b0000000101111010: out <= 16'h00AD;
			16'b0000000101111011: out <= 16'h00AC;
			16'b000000010111110x: out <= 16'h00AC;
			16'b000000010111111x: out <= 16'h00AB;
			16'b000000011000000x: out <= 16'h00AA;
			16'b000000011000001x: out <= 16'h00A9;
			16'b000000011000010x: out <= 16'h00A8;
			16'b0000000110000110: out <= 16'h00A8;
			16'b0000000110000111: out <= 16'h00A7;
			16'b0000000110001000: out <= 16'h00A7;
			16'b0000000110001001: out <= 16'h00A6;
			16'b0000000110001010: out <= 16'h00A6;
			16'b0000000110001011: out <= 16'h00A5;
			16'b000000011000110x: out <= 16'h00A5;
			16'b000000011000111x: out <= 16'h00A4;
			16'b000000011001000x: out <= 16'h00A3;
			16'b0000000110010010: out <= 16'h00A3;
			16'b0000000110010011: out <= 16'h00A2;
			16'b0000000110010100: out <= 16'h00A2;
			16'b0000000110010101: out <= 16'h00A1;
			16'b000000011001011x: out <= 16'h00A1;
			16'b000000011001100x: out <= 16'h00A0;
			16'b000000011001101x: out <= 16'h009F;
			16'b0000000110011100: out <= 16'h009F;
			16'b0000000110011101: out <= 16'h009E;
			16'b0000000110011110: out <= 16'h009E;
			16'b0000000110011111: out <= 16'h009D;
			16'b000000011010000x: out <= 16'h009D;
			16'b000000011010001x: out <= 16'h009C;
			16'b0000000110100100: out <= 16'h009C;
			16'b0000000110100101: out <= 16'h009B;
			16'b0000000110100110: out <= 16'h009B;
			16'b0000000110100111: out <= 16'h009A;
			16'b000000011010100x: out <= 16'h009A;
			16'b000000011010101x: out <= 16'h0099;
			16'b0000000110101100: out <= 16'h0099;
			16'b0000000110101101: out <= 16'h0098;
			16'b000000011010111x: out <= 16'h0098;
			16'b000000011011000x: out <= 16'h0097;
			16'b0000000110110010: out <= 16'h0097;
			16'b0000000110110011: out <= 16'h0096;
			16'b0000000110110100: out <= 16'h0096;
			16'b0000000110110101: out <= 16'h0095;
			16'b000000011011011x: out <= 16'h0095;
			16'b000000011011100x: out <= 16'h0094;
			16'b0000000110111010: out <= 16'h0094;
			16'b0000000110111011: out <= 16'h0093;
			16'b000000011011110x: out <= 16'h0093;
			16'b000000011011111x: out <= 16'h0092;
			16'b0000000111000000: out <= 16'h0092;
			16'b0000000111000001: out <= 16'h0091;
			16'b000000011100001x: out <= 16'h0091;
			16'b00000001110001xx: out <= 16'h0090;
			16'b000000011100100x: out <= 16'h008F;
			16'b0000000111001010: out <= 16'h008F;
			16'b0000000111001011: out <= 16'h008E;
			16'b000000011100110x: out <= 16'h008E;
			16'b000000011100111x: out <= 16'h008D;
			16'b0000000111010000: out <= 16'h008D;
			16'b0000000111010001: out <= 16'h008C;
			16'b000000011101001x: out <= 16'h008C;
			16'b0000000111010100: out <= 16'h008C;
			16'b0000000111010101: out <= 16'h008B;
			16'b000000011101011x: out <= 16'h008B;
			16'b000000011101100x: out <= 16'h008A;
			16'b0000000111011010: out <= 16'h008A;
			16'b0000000111011011: out <= 16'h0089;
			16'b000000011101110x: out <= 16'h0089;
			16'b0000000111011110: out <= 16'h0089;
			16'b0000000111011111: out <= 16'h0088;
			16'b000000011110000x: out <= 16'h0088;
			16'b000000011110001x: out <= 16'h0087;
			16'b000000011110010x: out <= 16'h0087;
			16'b000000011110011x: out <= 16'h0086;
			16'b000000011110100x: out <= 16'h0086;
			16'b000000011110101x: out <= 16'h0085;
			16'b0000000111101100: out <= 16'h0085;
			16'b0000000111101101: out <= 16'h0084;
			16'b000000011110111x: out <= 16'h0084;
			16'b0000000111110000: out <= 16'h0084;
			16'b0000000111110001: out <= 16'h0083;
			16'b000000011111001x: out <= 16'h0083;
			16'b0000000111110100: out <= 16'h0083;
			16'b0000000111110101: out <= 16'h0082;
			16'b000000011111011x: out <= 16'h0082;
			16'b0000000111111000: out <= 16'h0082;
			16'b0000000111111001: out <= 16'h0081;
			16'b000000011111101x: out <= 16'h0081;
			16'b0000000111111100: out <= 16'h0081;
			16'b0000000111111101: out <= 16'h0080;
			16'b000000011111111x: out <= 16'h0080;
			16'b0000001000000000: out <= 16'h0080;
			16'b0000001000000001: out <= 16'h007F;
			16'b000000100000001x: out <= 16'h007F;
			16'b0000001000000100: out <= 16'h007F;
			16'b0000001000000101: out <= 16'h007E;
			16'b000000100000011x: out <= 16'h007E;
			16'b0000001000001000: out <= 16'h007E;
			16'b0000001000001001: out <= 16'h007D;
			16'b000000100000101x: out <= 16'h007D;
			16'b0000001000001100: out <= 16'h007D;
			16'b0000001000001101: out <= 16'h007C;
			16'b000000100000111x: out <= 16'h007C;
			16'b0000001000010000: out <= 16'h007C;
			16'b0000001000010001: out <= 16'h007B;
			16'b000000100001001x: out <= 16'h007B;
			16'b0000001000010100: out <= 16'h007B;
			16'b0000001000010101: out <= 16'h007A;
			16'b000000100001011x: out <= 16'h007A;
			16'b000000100001100x: out <= 16'h007A;
			16'b000000100001101x: out <= 16'h0079;
			16'b000000100001110x: out <= 16'h0079;
			16'b000000100001111x: out <= 16'h0078;
			16'b000000100010000x: out <= 16'h0078;
			16'b0000001000100010: out <= 16'h0078;
			16'b0000001000100011: out <= 16'h0077;
			16'b000000100010010x: out <= 16'h0077;
			16'b0000001000100110: out <= 16'h0077;
			16'b0000001000100111: out <= 16'h0076;
			16'b00000010001010xx: out <= 16'h0076;
			16'b00000010001011xx: out <= 16'h0075;
			16'b000000100010111x: out <= 16'h0075;
			16'b0000001000110001: out <= 16'h0074;
			16'b000000100011001x: out <= 16'h0074;
			16'b0000001000110100: out <= 16'h0074;
			16'b0000001000110101: out <= 16'h0073;
			16'b000000100011011x: out <= 16'h0073;
			16'b000000100011100x: out <= 16'h0073;
			16'b000000100011101x: out <= 16'h0072;
			16'b000000100011110x: out <= 16'h0072;
			16'b0000001000111110: out <= 16'h0072;
			16'b0000001000111111: out <= 16'h0071;
			16'b00000010010000xx: out <= 16'h0071;
			16'b00000010010001xx: out <= 16'h0070;
			16'b000000100100100x: out <= 16'h0070;
			16'b000000100100101x: out <= 16'h006F;
			16'b000000100100110x: out <= 16'h006F;
			16'b0000001001001110: out <= 16'h006F;
			16'b0000001001001111: out <= 16'h006E;
			16'b00000010010100xx: out <= 16'h006E;
			16'b00000010010101xx: out <= 16'h006D;
			16'b000000100101100x: out <= 16'h006D;
			16'b000000100101101x: out <= 16'h006C;
			16'b000000100101110x: out <= 16'h006C;
			16'b0000001001011110: out <= 16'h006C;
			16'b0000001001011111: out <= 16'h006B;
			16'b00000010011000xx: out <= 16'h006B;
			16'b000000100110001x: out <= 16'h006B;
			16'b0000001001100101: out <= 16'h006A;
			16'b000000100110011x: out <= 16'h006A;
			16'b000000100110100x: out <= 16'h006A;
			16'b0000001001101010: out <= 16'h006A;
			16'b0000001001101011: out <= 16'h0069;
			16'b00000010011011xx: out <= 16'h0069;
			16'b000000100110111x: out <= 16'h0069;
			16'b0000001001110001: out <= 16'h0068;
			16'b000000100111001x: out <= 16'h0068;
			16'b000000100111010x: out <= 16'h0068;
			16'b0000001001110110: out <= 16'h0068;
			16'b0000001001110111: out <= 16'h0067;
			16'b00000010011110xx: out <= 16'h0067;
			16'b000000100111101x: out <= 16'h0067;
			16'b0000001001111101: out <= 16'h0066;
			16'b000000100111111x: out <= 16'h0066;
			16'b000000101000000x: out <= 16'h0066;
			16'b0000001010000010: out <= 16'h0066;
			16'b0000001010000011: out <= 16'h0065;
			16'b00000010100001xx: out <= 16'h0065;
			16'b000000101000011x: out <= 16'h0065;
			16'b0000001010001001: out <= 16'h0064;
			16'b000000101000101x: out <= 16'h0064;
			16'b00000010100011xx: out <= 16'h0064;
			16'b00000010100100xx: out <= 16'h0063;
			16'b000000101001010x: out <= 16'h0063;
			16'b000000101001011x: out <= 16'h0062;
			16'b00000010100110xx: out <= 16'h0062;
			16'b000000101001101x: out <= 16'h0062;
			16'b0000001010011101: out <= 16'h0061;
			16'b000000101001111x: out <= 16'h0061;
			16'b00000010101000xx: out <= 16'h0061;
			16'b00000010101001xx: out <= 16'h0060;
			16'b000000101010100x: out <= 16'h0060;
			16'b0000001010101010: out <= 16'h0060;
			16'b0000001010101011: out <= 16'h005F;
			16'b00000010101011xx: out <= 16'h005F;
			16'b000000101011000x: out <= 16'h005F;
			16'b000000101011001x: out <= 16'h005E;
			16'b00000010101101xx: out <= 16'h005E;
			16'b000000101011100x: out <= 16'h005E;
			16'b000000101011101x: out <= 16'h005D;
			16'b00000010101111xx: out <= 16'h005D;
			16'b000000101011111x: out <= 16'h005D;
			16'b0000001011000001: out <= 16'h005C;
			16'b000000101100001x: out <= 16'h005C;
			16'b00000010110001xx: out <= 16'h005C;
			16'b000000101100011x: out <= 16'h005C;
			16'b0000001011001001: out <= 16'h005B;
			16'b000000101100101x: out <= 16'h005B;
			16'b00000010110011xx: out <= 16'h005B;
			16'b000000101100111x: out <= 16'h005B;
			16'b0000001011010001: out <= 16'h005A;
			16'b000000101101001x: out <= 16'h005A;
			16'b00000010110101xx: out <= 16'h005A;
			16'b000000101101011x: out <= 16'h005A;
			16'b0000001011011001: out <= 16'h0059;
			16'b000000101101101x: out <= 16'h0059;
			16'b00000010110111xx: out <= 16'h0059;
			16'b000000101101111x: out <= 16'h0059;
			16'b0000001011100001: out <= 16'h0058;
			16'b000000101110001x: out <= 16'h0058;
			16'b00000010111001xx: out <= 16'h0058;
			16'b000000101110011x: out <= 16'h0058;
			16'b0000001011101001: out <= 16'h0057;
			16'b000000101110101x: out <= 16'h0057;
			16'b00000010111011xx: out <= 16'h0057;
			16'b000000101111000x: out <= 16'h0057;
			16'b000000101111001x: out <= 16'h0056;
			16'b00000010111101xx: out <= 16'h0056;
			16'b000000101111100x: out <= 16'h0056;
			16'b0000001011111010: out <= 16'h0056;
			16'b0000001011111011: out <= 16'h0055;
			16'b00000010111111xx: out <= 16'h0055;
			16'b00000011000000xx: out <= 16'h0055;
			16'b00000011000001xx: out <= 16'h0054;
			16'b00000011000010xx: out <= 16'h0054;
			16'b000000110000101x: out <= 16'h0054;
			16'b0000001100001101: out <= 16'h0053;
			16'b000000110000111x: out <= 16'h0053;
			16'b00000011000100xx: out <= 16'h0053;
			16'b000000110001010x: out <= 16'h0053;
			16'b000000110001011x: out <= 16'h0052;
			16'b0000001100011xxx: out <= 16'h0052;
			16'b0000001100100xxx: out <= 16'h0051;
			16'b00000011001001xx: out <= 16'h0051;
			16'b000000110010101x: out <= 16'h0050;
			16'b00000011001011xx: out <= 16'h0050;
			16'b00000011001100xx: out <= 16'h0050;
			16'b00000011001101xx: out <= 16'h004F;
			16'b00000011001110xx: out <= 16'h004F;
			16'b000000110011110x: out <= 16'h004F;
			16'b000000110011111x: out <= 16'h004E;
			16'b0000001101000xxx: out <= 16'h004E;
			16'b00000011010001xx: out <= 16'h004E;
			16'b0000001101001001: out <= 16'h004D;
			16'b000000110100101x: out <= 16'h004D;
			16'b00000011010011xx: out <= 16'h004D;
			16'b00000011010100xx: out <= 16'h004D;
			16'b00000011010101xx: out <= 16'h004C;
			16'b00000011010110xx: out <= 16'h004C;
			16'b000000110101110x: out <= 16'h004C;
			16'b0000001101011110: out <= 16'h004C;
			16'b0000001101011111: out <= 16'h004B;
			16'b0000001101100xxx: out <= 16'h004B;
			16'b00000011011001xx: out <= 16'h004B;
			16'b000000110110101x: out <= 16'h004A;
			16'b00000011011011xx: out <= 16'h004A;
			16'b00000011011100xx: out <= 16'h004A;
			16'b000000110111010x: out <= 16'h004A;
			16'b000000110111011x: out <= 16'h0049;
			16'b0000001101111xxx: out <= 16'h0049;
			16'b00000011011111xx: out <= 16'h0049;
			16'b000000111000001x: out <= 16'h0048;
			16'b00000011100001xx: out <= 16'h0048;
			16'b00000011100010xx: out <= 16'h0048;
			16'b000000111000110x: out <= 16'h0048;
			16'b0000001110001110: out <= 16'h0048;
			16'b0000001110001111: out <= 16'h0047;
			16'b0000001110010xxx: out <= 16'h0047;
			16'b00000011100110xx: out <= 16'h0047;
			16'b00000011100111xx: out <= 16'h0046;
			16'b0000001110100xxx: out <= 16'h0046;
			16'b00000011101001xx: out <= 16'h0046;
			16'b0000001110101001: out <= 16'h0045;
			16'b000000111010101x: out <= 16'h0045;
			16'b00000011101011xx: out <= 16'h0045;
			16'b00000011101100xx: out <= 16'h0045;
			16'b000000111011010x: out <= 16'h0045;
			16'b000000111011011x: out <= 16'h0044;
			16'b0000001110111xxx: out <= 16'h0044;
			16'b00000011110000xx: out <= 16'h0044;
			16'b00000011110001xx: out <= 16'h0043;
			16'b0000001111001xxx: out <= 16'h0043;
			16'b00000011110011xx: out <= 16'h0043;
			16'b000000111101000x: out <= 16'h0043;
			16'b0000001111010011: out <= 16'h0042;
			16'b00000011110101xx: out <= 16'h0042;
			16'b0000001111011xxx: out <= 16'h0042;
			16'b00000011110111xx: out <= 16'h0042;
			16'b0000001111100001: out <= 16'h0041;
			16'b000000111110001x: out <= 16'h0041;
			16'b00000011111001xx: out <= 16'h0041;
			16'b0000001111101xxx: out <= 16'h0041;
			16'b00000011111011xx: out <= 16'h0041;
			16'b0000001111110001: out <= 16'h0040;
			16'b000000111111001x: out <= 16'h0040;
			16'b00000011111101xx: out <= 16'h0040;
			16'b0000001111111xxx: out <= 16'h0040;
			16'b00000011111111xx: out <= 16'h0040;
			16'b0000010000000001: out <= 16'h003F;
			16'b000001000000001x: out <= 16'h003F;
			16'b00000100000001xx: out <= 16'h003F;
			16'b0000010000001xxx: out <= 16'h003F;
			16'b00000100000011xx: out <= 16'h003F;
			16'b0000010000010001: out <= 16'h003E;
			16'b000001000001001x: out <= 16'h003E;
			16'b00000100000101xx: out <= 16'h003E;
			16'b0000010000011xxx: out <= 16'h003E;
			16'b00000100000111xx: out <= 16'h003E;
			16'b000001000010001x: out <= 16'h003D;
			16'b00000100001001xx: out <= 16'h003D;
			16'b0000010000101xxx: out <= 16'h003D;
			16'b00000100001011xx: out <= 16'h003D;
			16'b000001000011000x: out <= 16'h003D;
			16'b0000010000110011: out <= 16'h003C;
			16'b00000100001101xx: out <= 16'h003C;
			16'b0000010000111xxx: out <= 16'h003C;
			16'b00000100010000xx: out <= 16'h003C;
			16'b000001000100001x: out <= 16'h003C;
			16'b0000010001000101: out <= 16'h003B;
			16'b000001000100011x: out <= 16'h003B;
			16'b0000010001001xxx: out <= 16'h003B;
			16'b00000100010100xx: out <= 16'h003B;
			16'b000001000101010x: out <= 16'h003B;
			16'b0000010001010110: out <= 16'h003B;
			16'b0000010001010111: out <= 16'h003A;
			16'b0000010001011xxx: out <= 16'h003A;
			16'b0000010001100xxx: out <= 16'h003A;
			16'b00000100011001xx: out <= 16'h003A;
			16'b000001000110101x: out <= 16'h0039;
			16'b00000100011011xx: out <= 16'h0039;
			16'b0000010001110xxx: out <= 16'h0039;
			16'b00000100011110xx: out <= 16'h0039;
			16'b000001000111110x: out <= 16'h0039;
			16'b000001000111111x: out <= 16'h0038;
			16'b000001001000xxxx: out <= 16'h0038;
			16'b0000010010001xxx: out <= 16'h0038;
			16'b00000100100011xx: out <= 16'h0038;
			16'b0000010010010011: out <= 16'h0037;
			16'b00000100100101xx: out <= 16'h0037;
			16'b0000010010011xxx: out <= 16'h0037;
			16'b0000010010100xxx: out <= 16'h0037;
			16'b0000010010101xxx: out <= 16'h0036;
			16'b0000010010110xxx: out <= 16'h0036;
			16'b00000100101110xx: out <= 16'h0036;
			16'b000001001011110x: out <= 16'h0036;
			16'b000001001011111x: out <= 16'h0035;
			16'b000001001100xxxx: out <= 16'h0035;
			16'b0000010011001xxx: out <= 16'h0035;
			16'b00000100110100xx: out <= 16'h0035;
			16'b0000010011010101: out <= 16'h0034;
			16'b000001001101011x: out <= 16'h0034;
			16'b0000010011011xxx: out <= 16'h0034;
			16'b0000010011100xxx: out <= 16'h0034;
			16'b00000100111010xx: out <= 16'h0034;
			16'b000001001110101x: out <= 16'h0034;
			16'b0000010011101101: out <= 16'h0033;
			16'b000001001110111x: out <= 16'h0033;
			16'b000001001111xxxx: out <= 16'h0033;
			16'b0000010011111xxx: out <= 16'h0033;
			16'b00000101000000xx: out <= 16'h0033;
			16'b000001010000011x: out <= 16'h0032;
			16'b0000010100001xxx: out <= 16'h0032;
			16'b0000010100010xxx: out <= 16'h0032;
			16'b00000101000110xx: out <= 16'h0032;
			16'b000001010001110x: out <= 16'h0032;
			16'b0000010100011110: out <= 16'h0032;
			16'b0000010100011111: out <= 16'h0031;
			16'b000001010010xxxx: out <= 16'h0031;
			16'b0000010100110xxx: out <= 16'h0031;
			16'b00000101001101xx: out <= 16'h0031;
			16'b000001010011101x: out <= 16'h0030;
			16'b00000101001111xx: out <= 16'h0030;
			16'b000001010100xxxx: out <= 16'h0030;
			16'b0000010101001xxx: out <= 16'h0030;
			16'b00000101010100xx: out <= 16'h0030;
			16'b000001010101011x: out <= 16'h002F;
			16'b0000010101011xxx: out <= 16'h002F;
			16'b000001010110xxxx: out <= 16'h002F;
			16'b0000010101101xxx: out <= 16'h002F;
			16'b00000101011011xx: out <= 16'h002F;
			16'b0000010101110011: out <= 16'h002E;
			16'b00000101011101xx: out <= 16'h002E;
			16'b0000010101111xxx: out <= 16'h002E;
			16'b000001011000xxxx: out <= 16'h002E;
			16'b0000010110001xxx: out <= 16'h002E;
			16'b0000010110010001: out <= 16'h002D;
			16'b000001011001001x: out <= 16'h002D;
			16'b00000101100101xx: out <= 16'h002D;
			16'b0000010110011xxx: out <= 16'h002D;
			16'b000001011010xxxx: out <= 16'h002D;
			16'b0000010110101xxx: out <= 16'h002D;
			16'b0000010110110001: out <= 16'h002C;
			16'b000001011011001x: out <= 16'h002C;
			16'b00000101101101xx: out <= 16'h002C;
			16'b0000010110111xxx: out <= 16'h002C;
			16'b000001011100xxxx: out <= 16'h002C;
			16'b0000010111001xxx: out <= 16'h002C;
			16'b000001011101001x: out <= 16'h002B;
			16'b00000101110101xx: out <= 16'h002B;
			16'b0000010111011xxx: out <= 16'h002B;
			16'b000001011110xxxx: out <= 16'h002B;
			16'b0000010111101xxx: out <= 16'h002B;
			16'b00000101111100xx: out <= 16'h002B;
			16'b0000010111110101: out <= 16'h002A;
			16'b000001011111011x: out <= 16'h002A;
			16'b0000010111111xxx: out <= 16'h002A;
			16'b000001100000xxxx: out <= 16'h002A;
			16'b0000011000010xxx: out <= 16'h002A;
			16'b00000110000101xx: out <= 16'h002A;
			16'b0000011000011001: out <= 16'h0029;
			16'b000001100001101x: out <= 16'h0029;
			16'b00000110000111xx: out <= 16'h0029;
			16'b000001100010xxxx: out <= 16'h0029;
			16'b0000011000110xxx: out <= 16'h0029;
			16'b00000110001110xx: out <= 16'h0029;
			16'b000001100011110x: out <= 16'h0029;
			16'b0000011000111110: out <= 16'h0029;
			16'b0000011000111111: out <= 16'h0028;
			16'b00000110010xxxxx: out <= 16'h0028;
			16'b000001100101xxxx: out <= 16'h0028;
			16'b0000011001011xxx: out <= 16'h0028;
			16'b00000110011000xx: out <= 16'h0028;
			16'b0000011001100111: out <= 16'h0027;
			16'b0000011001101xxx: out <= 16'h0027;
			16'b000001100111xxxx: out <= 16'h0027;
			16'b000001101000xxxx: out <= 16'h0027;
			16'b0000011010001xxx: out <= 16'h0027;
			16'b0000011010010001: out <= 16'h0026;
			16'b000001101001001x: out <= 16'h0026;
			16'b00000110100101xx: out <= 16'h0026;
			16'b0000011010011xxx: out <= 16'h0026;
			16'b000001101010xxxx: out <= 16'h0026;
			16'b0000011010110xxx: out <= 16'h0026;
			16'b00000110101110xx: out <= 16'h0026;
			16'b000001101011101x: out <= 16'h0026;
			16'b0000011010111101: out <= 16'h0025;
			16'b000001101011111x: out <= 16'h0025;
			16'b00000110110xxxxx: out <= 16'h0025;
			16'b000001101101xxxx: out <= 16'h0025;
			16'b0000011011100xxx: out <= 16'h0025;
			16'b00000110111011xx: out <= 16'h0024;
			16'b000001101111xxxx: out <= 16'h0024;
			16'b000001110000xxxx: out <= 16'h0024;
			16'b0000011100010xxx: out <= 16'h0024;
			16'b00000111000110xx: out <= 16'h0024;
			16'b000001110001101x: out <= 16'h0024;
			16'b0000011100011101: out <= 16'h0023;
			16'b000001110001111x: out <= 16'h0023;
			16'b00000111001xxxxx: out <= 16'h0023;
			16'b000001110100xxxx: out <= 16'h0023;
			16'b0000011101001xxx: out <= 16'h0023;
			16'b0000011101010001: out <= 16'h0022;
			16'b000001110101001x: out <= 16'h0022;
			16'b00000111010101xx: out <= 16'h0022;
			16'b0000011101011xxx: out <= 16'h0022;
			16'b00000111011xxxxx: out <= 16'h0022;
			16'b000001110111xxxx: out <= 16'h0022;
			16'b0000011110001xxx: out <= 16'h0021;
			16'b000001111001xxxx: out <= 16'h0021;
			16'b00000111101xxxxx: out <= 16'h0021;
			16'b000001111011xxxx: out <= 16'h0021;
			16'b000001111100001x: out <= 16'h0020;
			16'b00000111110001xx: out <= 16'h0020;
			16'b0000011111001xxx: out <= 16'h0020;
			16'b000001111101xxxx: out <= 16'h0020;
			16'b00000111111xxxxx: out <= 16'h0020;
			16'b000001111111xxxx: out <= 16'h0020;
			16'b0000100000000001: out <= 16'h001F;
			16'b000010000000001x: out <= 16'h001F;
			16'b00001000000001xx: out <= 16'h001F;
			16'b0000100000001xxx: out <= 16'h001F;
			16'b000010000001xxxx: out <= 16'h001F;
			16'b00001000001xxxxx: out <= 16'h001F;
			16'b000010000011xxxx: out <= 16'h001F;
			16'b0000100000111xxx: out <= 16'h001F;
			16'b0000100001000011: out <= 16'h001E;
			16'b00001000010001xx: out <= 16'h001E;
			16'b0000100001001xxx: out <= 16'h001E;
			16'b000010000101xxxx: out <= 16'h001E;
			16'b00001000011xxxxx: out <= 16'h001E;
			16'b000010000111xxxx: out <= 16'h001E;
			16'b0000100010000xxx: out <= 16'h001E;
			16'b0000100010001001: out <= 16'h001D;
			16'b000010001000101x: out <= 16'h001D;
			16'b00001000100011xx: out <= 16'h001D;
			16'b000010001001xxxx: out <= 16'h001D;
			16'b00001000101xxxxx: out <= 16'h001D;
			16'b000010001100xxxx: out <= 16'h001D;
			16'b0000100011001xxx: out <= 16'h001D;
			16'b00001000110101xx: out <= 16'h001C;
			16'b0000100011011xxx: out <= 16'h001C;
			16'b00001000111xxxxx: out <= 16'h001C;
			16'b00001001000xxxxx: out <= 16'h001C;
			16'b000010010001xxxx: out <= 16'h001C;
			16'b0000100100011xxx: out <= 16'h001C;
			16'b0000100100100101: out <= 16'h001B;
			16'b000010010010011x: out <= 16'h001B;
			16'b0000100100101xxx: out <= 16'h001B;
			16'b000010010011xxxx: out <= 16'h001B;
			16'b00001001010xxxxx: out <= 16'h001B;
			16'b000010010110xxxx: out <= 16'h001B;
			16'b0000100101110xxx: out <= 16'h001B;
			16'b00001001011110xx: out <= 16'h001B;
			16'b00001001011111xx: out <= 16'h001A;
			16'b0000100110xxxxxx: out <= 16'h001A;
			16'b00001001101xxxxx: out <= 16'h001A;
			16'b000010011100xxxx: out <= 16'h001A;
			16'b0000100111010xxx: out <= 16'h001A;
			16'b0000100111011001: out <= 16'h0019;
			16'b000010011101101x: out <= 16'h0019;
			16'b00001001110111xx: out <= 16'h0019;
			16'b00001001111xxxxx: out <= 16'h0019;
			16'b00001010000xxxxx: out <= 16'h0019;
			16'b000010100010xxxx: out <= 16'h0019;
			16'b0000101000110xxx: out <= 16'h0019;
			16'b00001010001110xx: out <= 16'h0019;
			16'b000010100011110x: out <= 16'h0019;
			16'b000010100011111x: out <= 16'h0018;
			16'b0000101001xxxxxx: out <= 16'h0018;
			16'b00001010100xxxxx: out <= 16'h0018;
			16'b000010101001xxxx: out <= 16'h0018;
			16'b0000101010100xxx: out <= 16'h0018;
			16'b00001010101001xx: out <= 16'h0018;
			16'b0000101010101011: out <= 16'h0017;
			16'b00001010101011xx: out <= 16'h0017;
			16'b000010101011xxxx: out <= 16'h0017;
			16'b0000101011xxxxxx: out <= 16'h0017;
			16'b00001011000xxxxx: out <= 16'h0017;
			16'b000010110001xxxx: out <= 16'h0017;
			16'b000010110010001x: out <= 16'h0016;
			16'b00001011001001xx: out <= 16'h0016;
			16'b0000101100101xxx: out <= 16'h0016;
			16'b000010110011xxxx: out <= 16'h0016;
			16'b0000101101xxxxxx: out <= 16'h0016;
			16'b00001011100xxxxx: out <= 16'h0016;
			16'b000010111001xxxx: out <= 16'h0016;
			16'b0000101110011xxx: out <= 16'h0016;
			16'b0000101110100011: out <= 16'h0015;
			16'b00001011101001xx: out <= 16'h0015;
			16'b0000101110101xxx: out <= 16'h0015;
			16'b000010111011xxxx: out <= 16'h0015;
			16'b0000101111xxxxxx: out <= 16'h0015;
			16'b00001100000xxxxx: out <= 16'h0015;
			16'b000011000010xxxx: out <= 16'h0015;
			16'b0000110000101xxx: out <= 16'h0015;
			16'b0000110000110001: out <= 16'h0014;
			16'b000011000011001x: out <= 16'h0014;
			16'b00001100001101xx: out <= 16'h0014;
			16'b0000110000111xxx: out <= 16'h0014;
			16'b0000110001xxxxxx: out <= 16'h0014;
			16'b0000110010xxxxxx: out <= 16'h0014;
			16'b00001100101xxxxx: out <= 16'h0014;
			16'b000011001011xxxx: out <= 16'h0014;
			16'b0000110011000xxx: out <= 16'h0014;
			16'b0000110011001101: out <= 16'h0013;
			16'b000011001100111x: out <= 16'h0013;
			16'b000011001101xxxx: out <= 16'h0013;
			16'b00001100111xxxxx: out <= 16'h0013;
			16'b0000110100xxxxxx: out <= 16'h0013;
			16'b00001101010xxxxx: out <= 16'h0013;
			16'b000011010110xxxx: out <= 16'h0013;
			16'b0000110101110xxx: out <= 16'h0013;
			16'b00001101011101xx: out <= 16'h0013;
			16'b000011010111101x: out <= 16'h0012;
			16'b00001101011111xx: out <= 16'h0012;
			16'b000011011xxxxxxx: out <= 16'h0012;
			16'b0000110111xxxxxx: out <= 16'h0012;
			16'b00001110000xxxxx: out <= 16'h0012;
			16'b000011100010xxxx: out <= 16'h0012;
			16'b0000111000110xxx: out <= 16'h0012;
			16'b0000111000111001: out <= 16'h0011;
			16'b000011100011101x: out <= 16'h0011;
			16'b00001110001111xx: out <= 16'h0011;
			16'b0000111001xxxxxx: out <= 16'h0011;
			16'b000011101xxxxxxx: out <= 16'h0011;
			16'b0000111011xxxxxx: out <= 16'h0011;
			16'b000011110001xxxx: out <= 16'h0010;
			16'b00001111001xxxxx: out <= 16'h0010;
			16'b000011111xxxxxxx: out <= 16'h0010;
			16'b0001000000000000: out <= 16'h0010;
			16'b0001000000000001: out <= 16'h000F;
			16'b000100000000001x: out <= 16'h000F;
			16'b00010000000001xx: out <= 16'h000F;
			16'b0001000000001xxx: out <= 16'h000F;
			16'b000100000001xxxx: out <= 16'h000F;
			16'b00010000001xxxxx: out <= 16'h000F;
			16'b0001000001xxxxxx: out <= 16'h000F;
			16'b000100001xxxxxxx: out <= 16'h000F;
			16'b000100010000xxxx: out <= 16'h000F;
			16'b000100010001000x: out <= 16'h000F;
			16'b000100010001001x: out <= 16'h000E;
			16'b00010001000101xx: out <= 16'h000E;
			16'b0001000100011xxx: out <= 16'h000E;
			16'b00010001001xxxxx: out <= 16'h000E;
			16'b0001000101xxxxxx: out <= 16'h000E;
			16'b000100011xxxxxxx: out <= 16'h000E;
			16'b0001000xxxxxxxxx: out <= 16'h000E;
			16'b0001001000xxxxxx: out <= 16'h000E;
			16'b0001001001000xxx: out <= 16'h000E;
			16'b000100100100100x: out <= 16'h000E;
			16'b000100100100101x: out <= 16'h000D;
			16'b00010010010011xx: out <= 16'h000D;
			16'b000100100101xxxx: out <= 16'h000D;
			16'b00010010011xxxxx: out <= 16'h000D;
			16'b000100101xxxxxxx: out <= 16'h000D;
			16'b000100110xxxxxxx: out <= 16'h000D;
			16'b00010011100xxxxx: out <= 16'h000D;
			16'b000100111010xxxx: out <= 16'h000D;
			16'b000100111011000x: out <= 16'h000D;
			16'b000100111011001x: out <= 16'h000C;
			16'b00010011101101xx: out <= 16'h000C;
			16'b0001001110111xxx: out <= 16'h000C;
			16'b0001001111xxxxxx: out <= 16'h000C;
			16'b00010100xxxxxxxx: out <= 16'h000C;
			16'b0001010100xxxxxx: out <= 16'h000C;
			16'b000101010100xxxx: out <= 16'h000C;
			16'b00010101010100xx: out <= 16'h000C;
			16'b000101010101010x: out <= 16'h000C;
			16'b000101010101011x: out <= 16'h000B;
			16'b0001010101011xxx: out <= 16'h000B;
			16'b00010101011xxxxx: out <= 16'h000B;
			16'b000101011xxxxxxx: out <= 16'h000B;
			16'b00010110xxxxxxxx: out <= 16'h000B;
			16'b0001011100xxxxxx: out <= 16'h000B;
			16'b00010111010000xx: out <= 16'h000B;
			16'b000101110100010x: out <= 16'h000B;
			16'b000101110100011x: out <= 16'h000A;
			16'b0001011101001xxx: out <= 16'h000A;
			16'b000101110101xxxx: out <= 16'h000A;
			16'b00010111011xxxxx: out <= 16'h000A;
			16'b000101111xxxxxxx: out <= 16'h000A;
			16'b00011000xxxxxxxx: out <= 16'h000A;
			16'b000110010xxxxxxx: out <= 16'h000A;
			16'b000110011000xxxx: out <= 16'h000A;
			16'b0001100110010xxx: out <= 16'h000A;
			16'b000110011001100x: out <= 16'h000A;
			16'b000110011001101x: out <= 16'h0009;
			16'b00011001100111xx: out <= 16'h0009;
			16'b00011001101xxxxx: out <= 16'h0009;
			16'b0001100111xxxxxx: out <= 16'h0009;
			16'b0001101xxxxxxxxx: out <= 16'h0009;
			16'b0001110000xxxxxx: out <= 16'h0009;
			16'b00011100010xxxxx: out <= 16'h0009;
			16'b000111000110xxxx: out <= 16'h0009;
			16'b000111000111000x: out <= 16'h0009;
			16'b000111000111001x: out <= 16'h0008;
			16'b00011100011101xx: out <= 16'h0008;
			16'b0001110001111xxx: out <= 16'h0008;
			16'b000111001xxxxxxx: out <= 16'h0008;
			16'b00011101xxxxxxxx: out <= 16'h0008;
			16'b0001111xxxxxxxxx: out <= 16'h0008;
			16'b0010000000000000: out <= 16'h0008;
			16'b0010000000000001: out <= 16'h0007;
			16'b001000000000001x: out <= 16'h0007;
			16'b00100000000001xx: out <= 16'h0007;
			16'b0010000000001xxx: out <= 16'h0007;
			16'b001000000001xxxx: out <= 16'h0007;
			16'b00100000001xxxxx: out <= 16'h0007;
			16'b0010000001xxxxxx: out <= 16'h0007;
			16'b001000001xxxxxxx: out <= 16'h0007;
			16'b00100001xxxxxxxx: out <= 16'h0007;
			16'b0010001xxxxxxxxx: out <= 16'h0007;
			16'b001001000xxxxxxx: out <= 16'h0007;
			16'b001001001000xxxx: out <= 16'h0007;
			16'b001001001001000x: out <= 16'h0007;
			16'b0010010010010010: out <= 16'h0007;
			16'b0010010010010011: out <= 16'h0006;
			16'b00100100100101xx: out <= 16'h0006;
			16'b0010010010011xxx: out <= 16'h0006;
			16'b00100100101xxxxx: out <= 16'h0006;
			16'b0010010011xxxxxx: out <= 16'h0006;
			16'b00100101xxxxxxxx: out <= 16'h0006;
			16'b0010011xxxxxxxxx: out <= 16'h0006;
			16'b0010100xxxxxxxxx: out <= 16'h0006;
			16'b001010100xxxxxxx: out <= 16'h0006;
			16'b00101010100xxxxx: out <= 16'h0006;
			16'b0010101010100xxx: out <= 16'h0006;
			16'b001010101010100x: out <= 16'h0006;
			16'b0010101010101010: out <= 16'h0006;
			16'b0010101010101011: out <= 16'h0005;
			16'b00101010101011xx: out <= 16'h0005;
			16'b001010101011xxxx: out <= 16'h0005;
			16'b0010101011xxxxxx: out <= 16'h0005;
			16'b00101011xxxxxxxx: out <= 16'h0005;
			16'b001011xxxxxxxxxx: out <= 16'h0005;
			16'b0011000xxxxxxxxx: out <= 16'h0005;
			16'b00110010xxxxxxxx: out <= 16'h0005;
			16'b00110011000xxxxx: out <= 16'h0005;
			16'b001100110010xxxx: out <= 16'h0005;
			16'b00110011001100xx: out <= 16'h0005;
			16'b00110011001101xx: out <= 16'h0004;
			16'b0011001100111xxx: out <= 16'h0004;
			16'b0011001101xxxxxx: out <= 16'h0004;
			16'b001100111xxxxxxx: out <= 16'h0004;
			16'b001101xxxxxxxxxx: out <= 16'h0004;
			16'b00111xxxxxxxxxxx: out <= 16'h0004;
			16'b0100000000000000: out <= 16'h0004;
			16'b0100000000000001: out <= 16'h0003;
			16'b010000000000001x: out <= 16'h0003;
			16'b010000000000001x: out <= 16'h0003;
			16'b01000000000001xx: out <= 16'h0003;
			16'b0100000000001xxx: out <= 16'h0003;
			16'b010000000001xxxx: out <= 16'h0003;
			16'b01000000001xxxxx: out <= 16'h0003;
			16'b0100000001xxxxxx: out <= 16'h0003;
			16'b010000001xxxxxxx: out <= 16'h0003;
			16'b01000001xxxxxxxx: out <= 16'h0003;
			16'b0100001xxxxxxxxx: out <= 16'h0003;
			16'b010001xxxxxxxxxx: out <= 16'h0003;
			16'b01001xxxxxxxxxxx: out <= 16'h0003;
			16'b010100xxxxxxxxxx: out <= 16'h0003;
			16'b01010100xxxxxxxx: out <= 16'h0003;
			16'b0101010100xxxxxx: out <= 16'h0003;
			16'b010101010100xxxx: out <= 16'h0003;
			16'b01010101010100xx: out <= 16'h0003;
			16'b010101010101010x: out <= 16'h0003;
			16'b010101010101011x: out <= 16'h0002;
			16'b010101010101011x: out <= 16'h0002;
			16'b0101010101011xxx: out <= 16'h0002;
			16'b01010101011xxxxx: out <= 16'h0002;
			16'b010101011xxxxxxx: out <= 16'h0002;
			16'b0101011xxxxxxxxx: out <= 16'h0002;
			16'b01011xxxxxxxxxxx: out <= 16'h0002;
			16'b011xxxxxxxxxxxxx: out <= 16'h0002;
			16'b1000000000000000: out <= 16'h0002;
			16'b1000000000000001: out <= 16'h0001;
			16'b100000000000001x: out <= 16'h0001;
			16'b10000000000001xx: out <= 16'h0001;
			16'b1000000000001xxx: out <= 16'h0001;
			16'b100000000001xxxx: out <= 16'h0001;
			16'b10000000001xxxxx: out <= 16'h0001;
			16'b1000000001xxxxxx: out <= 16'h0001;
			16'b100000001xxxxxxx: out <= 16'h0001;
			16'b10000001xxxxxxxx: out <= 16'h0001;
			16'b1000001xxxxxxxxx: out <= 16'h0001;
			16'b100001xxxxxxxxxx: out <= 16'h0001;
			16'b10001xxxxxxxxxxx: out <= 16'h0001;
			16'b1001xxxxxxxxxxxx: out <= 16'h0001;
			16'b101xxxxxxxxxxxxx: out <= 16'h0001;
			16'b11xxxxxxxxxxxxxx: out <= 16'h0001;
			default: out <= 16'h0000;
		endcase
	end
	
	always @ (posedge clk)
	begin
		if (en)
		begin
			if (a == b)
				xyouti <= 32'h10000;
			else if (b == 16'h0001)
				xyouti <= { a, 16'h0000 };
			else
				xyouti <= temp;
		end
		xyout <= xyouti;
	end
	
endmodule

module mult (
	input wire [15:0] a,
	input wire [15:0] b,
	output reg [31:0] result
	);
	
	integer i;
	
	always @ (a or b)
	begin
		result = 0;
		for (i = 0; i < 16; i = i + 1) // 이게 합성이 되나??
		if (a[i] == 1'b1)
			result = result + ( b << i );
	end
	
endmodule
